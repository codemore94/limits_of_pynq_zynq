module Transformer(
		   input clk,
		   input rst,
		   input reg[DATA_WIDTH-1:0],
		   output reg[DATA_WIDTH-1:0]
);

   reg					     attention_out[DATA_WIDTH-1:0];
   reg					     ff_out[DATA_WIDTH-1:0];
   reg					     norm_out[DATA_WIDTH-1:0];
end module;
   
   
   
   
